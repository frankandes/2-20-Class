type carry_array is array(N-1 downto 1) of std_logic_vector(N-1 downto 0);
type and_array is array(N-1 downto 0) of std_logic_vector(N-1 downto 0);
.
.
.
a : and_array
.
.
.
begin